Start Writing Synthesis Report
---------------------------------------------------------------------------------

DSP Final Report (the ' indicates corresponding REG is set)
+--------------+--------------+--------+--------+--------+--------+--------+------+------+------+------+-------+------+------+
|Module Name   | DSP Mapping  | A Size | B Size | C Size | D Size | P Size | AREG | BREG | CREG | DREG | ADREG | MREG | PREG | 
+--------------+--------------+--------+--------+--------+--------+--------+------+------+------+------+-------+------+------+
|fp_multiplier | A*B          | 24     | 17     | -      | -      | 48     | 0    | 0    | -    | -    | -     | 0    | 0    | 
|fp_multiplier | PCIN>>17+A*B | 0      | 7      | -      | -      | 31     | 0    | 0    | -    | -    | -     | 0    | 0    | 
+--------------+--------------+--------+--------+--------+--------+--------+------+------+------+------+-------+------+------+


Report BlackBoxes: 
+-+--------------+----------+
| |BlackBox name |Instances |
+-+--------------+----------+
+-+--------------+----------+

Report Cell Usage: 
+------+--------+------+
|      |Cell    |Count |
+------+--------+------+
|1     |CARRY4  |     2|
|2     |DSP48E1 |     2|
|3     |LUT2    |     5|
|4     |LUT3    |    26|
|5     |LUT4    |     6|
|6     |LUT5    |     1|
|7     |IBUF    |    64|
|8     |OBUF    |    32|
+------+--------+------+

Report Instance Areas: 
+------+---------+-------+------+
|      |Instance |Module |Cells |
+------+---------+-------+------+
|1     |top      |       |   138|
+------+---------+-------+------+
---------------------------------------------------------------------------------
Finished Writing Synthesis Report

